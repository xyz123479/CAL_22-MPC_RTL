module TRANSFORMER #(
  parameter[0:7]   ROOT_IDX = 8'd21,
  parameter[0:255] BASE_IDX = {
    8'd11, 8'd11, 8'd23, 8'd11, 8'd07, 8'd07, 8'd07, 8'd15,
    8'd11, 8'd11, 8'd07, 8'd19, 8'd15, 8'd15, 8'd23, 8'd23,
    8'd19, 8'd19, 8'd23, 8'd23, 8'd23, 8'd21, 8'd23, 8'd21,
    8'd27, 8'd27, 8'd23, 8'd19, 8'd31, 8'd11, 8'd23, 8'd23
  },
  parameter[0:255] SHIFT_VAL = {
    8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,
    8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,
    8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,
    8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0,  8'd0
  },
  parameter[0:2047] SCAN_ROW = {
    8'd4, 8'd4, 8'd4, 8'd2, 8'd4, 8'd3, 8'd3, 8'd3,
    8'd4, 8'd2, 8'd2, 8'd2, 8'd2, 8'd2, 8'd2, 8'd4,
    8'd3, 8'd3, 8'd3, 8'd4, 8'd3, 8'd5, 8'd5, 8'd5,
    8'd5, 8'd5, 8'd5, 8'd5, 8'd6, 8'd6, 8'd6, 8'd6,
    8'd6, 8'd6, 8'd6, 8'd7, 8'd7, 8'd7, 8'd7, 8'd7,
    8'd7, 8'd7, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd0,
    8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd0,
    8'd1, 8'd1, 8'd1, 8'd0, 8'd1, 8'd1, 8'd1, 8'd1,
    8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0,
    8'd5, 8'd5, 8'd3, 8'd5, 8'd5, 8'd5, 8'd5, 8'd2,
    8'd7, 8'd4, 8'd7, 8'd4, 8'd6, 8'd6, 8'd4, 8'd5,
    8'd1, 8'd0, 8'd0, 8'd0, 8'd7, 8'd6, 8'd7, 8'd7,
    8'd4, 8'd5, 8'd5, 8'd7, 8'd2, 8'd7, 8'd7, 8'd7,
    8'd4, 8'd3, 8'd5, 8'd3, 8'd6, 8'd6, 8'd6, 8'd6,
    8'd6, 8'd5, 8'd2, 8'd2, 8'd4, 8'd4, 8'd4, 8'd7,
    8'd7, 8'd3, 8'd5, 8'd6, 8'd6, 8'd6, 8'd5, 8'd6,
    8'd6, 8'd5, 8'd0, 8'd0, 8'd0, 8'd1, 8'd0, 8'd0,
    8'd2, 8'd2, 8'd2, 8'd2, 8'd4, 8'd5, 8'd5, 8'd4,
    8'd2, 8'd3, 8'd0, 8'd0, 8'd4, 8'd2, 8'd2, 8'd0,
    8'd0, 8'd4, 8'd4, 8'd4, 8'd4, 8'd3, 8'd4, 8'd4,
    8'd4, 8'd3, 8'd3, 8'd2, 8'd4, 8'd7, 8'd3, 8'd0,
    8'd0, 8'd0, 8'd2, 8'd4, 8'd1, 8'd1, 8'd2, 8'd0,
    8'd1, 8'd1, 8'd1, 8'd3, 8'd7, 8'd6, 8'd6, 8'd6,
    8'd7, 8'd4, 8'd3, 8'd3, 8'd5, 8'd2, 8'd3, 8'd3,
    8'd6, 8'd5, 8'd5, 8'd3, 8'd5, 8'd7, 8'd5, 8'd4,
    8'd3, 8'd2, 8'd6, 8'd5, 8'd5, 8'd2, 8'd3, 8'd7,
    8'd3, 8'd6, 8'd2, 8'd3, 8'd3, 8'd3, 8'd6, 8'd2,
    8'd2, 8'd4, 8'd7, 8'd6, 8'd6, 8'd6, 8'd2, 8'd2,
    8'd2, 8'd5, 8'd4, 8'd2, 8'd3, 8'd3, 8'd2, 8'd7,
    8'd7, 8'd7, 8'd7, 8'd6, 8'd6, 8'd5, 8'd3, 8'd3,
    8'd7, 8'd7, 8'd7, 8'd7, 8'd1, 8'd1, 8'd1, 8'd4,
    8'd1, 8'd1, 8'd1, 8'd1, 8'd1, 8'd1, 8'd1, 8'd1
  },
  parameter[0:2047] SCAN_COL = {
    8'd31, 8'd27, 8'd04, 8'd20, 8'd08, 8'd27, 8'd12, 8'd04,
    8'd12, 8'd27, 8'd08, 8'd16, 8'd04, 8'd12, 8'd31, 8'd16,
    8'd16, 8'd08, 8'd31, 8'd20, 8'd20, 8'd20, 8'd31, 8'd27,
    8'd12, 8'd08, 8'd16, 8'd04, 8'd20, 8'd31, 8'd16, 8'd08,
    8'd27, 8'd12, 8'd04, 8'd04, 8'd20, 8'd16, 8'd31, 8'd08,
    8'd27, 8'd12, 8'd16, 8'd16, 8'd08, 8'd08, 8'd12, 8'd12,
    8'd27, 8'd27, 8'd31, 8'd31, 8'd04, 8'd04, 8'd20, 8'd20,
    8'd17, 8'd21, 8'd09, 8'd00, 8'd00, 8'd05, 8'd13, 8'd24,
    8'd07, 8'd11, 8'd22, 8'd26, 8'd30, 8'd15, 8'd19, 8'd03,
    8'd13, 8'd21, 8'd00, 8'd28, 8'd17, 8'd01, 8'd05, 8'd00,
    8'd07, 8'd06, 8'd15, 8'd00, 8'd23, 8'd00, 8'd23, 8'd15,
    8'd28, 8'd28, 8'd05, 8'd06, 8'd06, 8'd14, 8'd22, 8'd10,
    8'd25, 8'd24, 8'd09, 8'd25, 8'd24, 8'd29, 8'd14, 8'd30,
    8'd14, 8'd23, 8'd22, 8'd14, 8'd13, 8'd28, 8'd21, 8'd05,
    8'd06, 8'd07, 8'd07, 8'd03, 8'd02, 8'd18, 8'd10, 8'd18,
    8'd02, 8'd06, 8'd30, 8'd29, 8'd26, 8'd11, 8'd18, 8'd19,
    8'd03, 8'd25, 8'd02, 8'd10, 8'd01, 8'd01, 8'd09, 8'd29,
    8'd22, 8'd19, 8'd15, 8'd11, 8'd11, 8'd10, 8'd02, 8'd03,
    8'd17, 8'd29, 8'd18, 8'd17, 8'd26, 8'd26, 8'd30, 8'd14,
    8'd13, 8'd17, 8'd24, 8'd09, 8'd01, 8'd01, 8'd05, 8'd21,
    8'd28, 8'd28, 8'd17, 8'd25, 8'd29, 8'd03, 8'd25, 8'd21,
    8'd25, 8'd24, 8'd09, 8'd19, 8'd10, 8'd02, 8'd01, 8'd23,
    8'd23, 8'd14, 8'd25, 8'd18, 8'd19, 8'd10, 8'd01, 8'd17,
    8'd11, 8'd13, 8'd13, 8'd21, 8'd14, 8'd28, 8'd24, 8'd05,
    8'd25, 8'd03, 8'd19, 8'd03, 8'd23, 8'd00, 8'd00, 8'd15,
    8'd09, 8'd18, 8'd18, 8'd26, 8'd29, 8'd29, 8'd02, 8'd26,
    8'd10, 8'd02, 8'd02, 8'd11, 8'd19, 8'd22, 8'd07, 8'd05,
    8'd21, 8'd22, 8'd23, 8'd22, 8'd30, 8'd15, 8'd14, 8'd23,
    8'd10, 8'd06, 8'd07, 8'd06, 8'd07, 8'd15, 8'd13, 8'd13,
    8'd28, 8'd21, 8'd05, 8'd24, 8'd09, 8'd11, 8'd26, 8'd30,
    8'd24, 8'd01, 8'd09, 8'd17, 8'd29, 8'd06, 8'd18, 8'd30,
    8'd03, 8'd07, 8'd11, 8'd26, 8'd22, 8'd30, 8'd15, 8'd19
  }
) (
  input [255:0] data_i,

  output [255:0] data_o
);
// synopsys template

  wire [  7:0] root;
  wire [247:0] data;
  wire [247:0] pred;
  PREDICTOR #(
    .ROOT_IDX  (ROOT_IDX),
    .BASE_IDX  (BASE_IDX),
    .SHIFT_VAL (SHIFT_VAL)
  ) PRED0 (
    .data_i	(data_i),
    .root_o	(root),
    .data_o (data),
    .pred_o (pred)
  );

  wire [247:0] diff_o;
  SUBTRACTOR SUB0 (
    .data_i (data),
    .pred_i (pred),
    .diff_o (diff_o)
  );

  wire [255:0] diff_i;
  wire [255:0] bpx;
  assign diff_i = { root, diff_o };
  DBX DBX0 (
    .diff_i (diff_i),
    .bpx_o	(bpx)
  );

  wire [255:0] scanned;
  SCAN #(
   .SCAN_COL (SCAN_COL),
   .SCAN_ROW (SCAN_ROW)
  ) SCAN0 (
    .bpx_i		(bpx),
    .scanned_o(scanned)
  );

  assign data_o = scanned;

endmodule


